module yAlu(z, ex, a, b, op);
input [31:0] a, b;
input [2:0] op;
output [31:0] z;
output ex;
wire [31:0] a0, a1, a2, slt;
wire [15:0] z16;
wire [7:0] z8;
wire [3:0] z4;
wire [1:0] z2;
wire z1;
assign slt[31:1] = 0; // not supported
//assign ex = 0;// not supported

yArith cal[31:0](a2, cout, a, b, op[2]);
and Alu_and[31:0](a0, a, b);
or Alu_or[31:0](a1, a, b);

xor Alu_xor(xoro, a[31], b[31]);
yMux1 Alu_slt(slt[0],a[31], a2[31], xoro);

yMux4to1 #(32) select(z, a0, a1, a2, slt, op[1:0]); 

or or16[15:0](z16, z[15:0], z[31:16]);
or or8[7:0](z8, z16[7:0], z16[15:8]);
or or4[3:0](z4, z8[3:0], z8[7:4]);
or or2[1:0](z2, z4[1:0], z4[3:2]);
or or1(z1, z2[1], z2[0]);
not mynot(ex, z2);
 
endmodule